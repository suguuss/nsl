library ieee;
use ieee.std_logic_1164.all;

library nsl_cuff, nsl_line_coding, nsl_io;
use nsl_cuff.protocol.all;

entity cuff_receiver is
    generic (
        lane_count_c           : natural;
        input_fixed_delay_ps_c : natural := 0;
        has_input_alignment_c  : boolean := true;
        sdr_ddr_c              : string  := "ddr"
    );
    port (
        clock_i         : in std_ulogic;
        gearbox_clock_i : in std_ulogic := '0';
        bit_clock_i     : in std_ulogic;
        reset_n_i       : in std_ulogic;

        serdes_strobe_i : in std_ulogic := '0';

        pad_i  : in  std_ulogic_vector(0 to lane_count_c - 1);
        lane_o : out cuff_code_vector(0 to lane_count_c - 1);

        align_restart_i : in  std_ulogic;
        align_valid_i   : in  std_ulogic_vector(0 to lane_count_c - 1);
        align_ready_o   : out std_ulogic_vector(0 to lane_count_c - 1)
    );
end entity;

architecture xc6 of cuff_receiver is
    component input_delay_variable is
        port (
            clock_i     : in  std_ulogic;
            bit_clock_i : in  std_ulogic;
            reset_n_i   : in  std_ulogic;
            mark_o      : out std_ulogic;
            shift_i     : in  std_ulogic;

            data_i : in  std_ulogic;
            data_o : out std_ulogic
        );
    end component;
begin

    iter : for i in 0 to lane_count_c - 1
        generate
        signal delayed_s, delay_shift_s, delay_mark_s, slip_shift_s, slip_mark_s : std_ulogic;
    begin
        with_aligner : if has_input_alignment_c
            generate
            aligner : nsl_io.delay.input_delay_aligner
            generic map(
                stabilization_delay_c => 7,
                stabilization_cycle_c => 6
            )
            port map(
                clock_i   => gearbox_clock_i,
                reset_n_i => reset_n_i,

                delay_shift_o  => delay_shift_s,
                delay_mark_i   => delay_mark_s,
                serdes_shift_o => slip_shift_s,
                serdes_mark_i  => slip_mark_s,

                restart_i => align_restart_i,
                valid_i   => align_valid_i(i),
                ready_o   => align_ready_o(i)
            );

            -- delayer : nsl_io.delay.input_delay_variable
            xc6_delayer : input_delay_variable
            port map(
                clock_i     => gearbox_clock_i,
                reset_n_i   => reset_n_i,
                bit_clock_i => bit_clock_i,
                mark_o      => delay_mark_s,
                shift_i     => delay_shift_s,
                data_i      => pad_i(i),
                data_o      => delayed_s
            );
        end generate;

        without_aligner : if not has_input_alignment_c
            generate
            delay : nsl_io.delay.input_delay_fixed
            generic map(
                delay_ps_c => input_fixed_delay_ps_c,
                is_ddr_c   => true
            )
            port map(
                data_i => pad_i(i),
                data_o => delayed_s
            );

            align_ready_o(i) <= '1';
        end generate;

        ddr_gen : if sdr_ddr_c = "ddr" generate
            deserializer : nsl_io.serdes.serdes_ddr10_input
            port map(
                word_clock_i => clock_i,
                bit_clock_i  => bit_clock_i,
                reset_n_i    => reset_n_i,
                parallel_o   => lane_o(i),
                serial_i     => delayed_s,
                bitslip_i    => slip_shift_s,
                mark_o       => slip_mark_s
            );
        end generate;

        sdr_gen : if sdr_ddr_c = "sdr" generate
            deserializer : nsl_io.serdes.serdes_sdr10_input
            port map(
                word_clock_i    => clock_i,
                gearbox_clock_i => gearbox_clock_i,
                bit_clock_i     => bit_clock_i,
                reset_n_i       => reset_n_i,
                serdes_strobe_i => serdes_strobe_i,
                parallel_o      => lane_o(i),
                serial_i        => delayed_s,
                bitslip_i       => slip_shift_s,
                mark_o          => slip_mark_s
            );
        end generate;
    end generate;

end architecture;
